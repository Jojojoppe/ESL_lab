// nios.v

// Generated using ACDS version 13.1 162 at 2021.06.22.13:12:26

`timescale 1 ps / 1 ps
module nios (
		input  wire       clk_clk,                        //                        clk.clk
		input  wire       reset_reset_n,                  //                      reset.reset_n
		input  wire       uart_0_external_connection_rxd, // uart_0_external_connection.rxd
		output wire       uart_0_external_connection_txd, //                           .txd
		input  wire       enc1a_encoder_a,                //                      enc1a.encoder_a
		input  wire       enc1b_encoder_b,                //                      enc1b.encoder_b
		input  wire       enc2a_encoder_a,                //                      enc2a.encoder_a
		input  wire       enc2b_encoder_b,                //                      enc2b.encoder_b
		output wire [7:0] enc1leds_leds,                  //                   enc1leds.leds
		output wire [7:0] enc2leds_leds,                  //                   enc2leds.leds
		inout  wire       pwma_ina,                       //                       pwma.ina
		inout  wire       pwma_inb,                       //                           .inb
		output wire       pwma_inc,                       //                           .inc
		inout  wire       pwmb_ina,                       //                       pwmb.ina
		inout  wire       pwmb_inb,                       //                           .inb
		output wire       pwmb_inc                        //                           .inc
	);

	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_esl_pwm_0_s0_writedata;                     // mm_interconnect_0:esl_pwm_0_s0_writedata -> esl_pwm_0:slave_writedata
	wire   [7:0] mm_interconnect_0_esl_pwm_0_s0_address;                       // mm_interconnect_0:esl_pwm_0_s0_address -> esl_pwm_0:slave_address
	wire         mm_interconnect_0_esl_pwm_0_s0_write;                         // mm_interconnect_0:esl_pwm_0_s0_write -> esl_pwm_0:slave_write
	wire         mm_interconnect_0_esl_pwm_0_s0_read;                          // mm_interconnect_0:esl_pwm_0_s0_read -> esl_pwm_0:slave_read
	wire  [31:0] mm_interconnect_0_esl_pwm_0_s0_readdata;                      // esl_pwm_0:slave_readdata -> mm_interconnect_0:esl_pwm_0_s0_readdata
	wire   [3:0] mm_interconnect_0_esl_pwm_0_s0_byteenable;                    // mm_interconnect_0:esl_pwm_0_s0_byteenable -> esl_pwm_0:slave_byteenable
	wire  [31:0] mm_interconnect_0_esl_pwm_1_s0_writedata;                     // mm_interconnect_0:esl_pwm_1_s0_writedata -> esl_pwm_1:slave_writedata
	wire   [7:0] mm_interconnect_0_esl_pwm_1_s0_address;                       // mm_interconnect_0:esl_pwm_1_s0_address -> esl_pwm_1:slave_address
	wire         mm_interconnect_0_esl_pwm_1_s0_write;                         // mm_interconnect_0:esl_pwm_1_s0_write -> esl_pwm_1:slave_write
	wire         mm_interconnect_0_esl_pwm_1_s0_read;                          // mm_interconnect_0:esl_pwm_1_s0_read -> esl_pwm_1:slave_read
	wire  [31:0] mm_interconnect_0_esl_pwm_1_s0_readdata;                      // esl_pwm_1:slave_readdata -> mm_interconnect_0:esl_pwm_1_s0_readdata
	wire   [3:0] mm_interconnect_0_esl_pwm_1_s0_byteenable;                    // mm_interconnect_0:esl_pwm_1_s0_byteenable -> esl_pwm_1:slave_byteenable
	wire  [31:0] mm_interconnect_0_esl_encoder_0_s0_writedata;                 // mm_interconnect_0:esl_encoder_0_s0_writedata -> esl_encoder_0:slave_writedata
	wire   [7:0] mm_interconnect_0_esl_encoder_0_s0_address;                   // mm_interconnect_0:esl_encoder_0_s0_address -> esl_encoder_0:slave_address
	wire         mm_interconnect_0_esl_encoder_0_s0_write;                     // mm_interconnect_0:esl_encoder_0_s0_write -> esl_encoder_0:slave_write
	wire         mm_interconnect_0_esl_encoder_0_s0_read;                      // mm_interconnect_0:esl_encoder_0_s0_read -> esl_encoder_0:slave_read
	wire  [31:0] mm_interconnect_0_esl_encoder_0_s0_readdata;                  // esl_encoder_0:slave_readdata -> mm_interconnect_0:esl_encoder_0_s0_readdata
	wire   [3:0] mm_interconnect_0_esl_encoder_0_s0_byteenable;                // mm_interconnect_0:esl_encoder_0_s0_byteenable -> esl_encoder_0:slave_byteenable
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                       // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                         // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                      // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                           // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                        // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [16:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_readdatavalid;                // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [16:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                        // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                          // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_chipselect;                       // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire         mm_interconnect_0_uart_0_s1_write;                            // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire         mm_interconnect_0_uart_0_s1_read;                             // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                         // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                    // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;         // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;        // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire  [31:0] mm_interconnect_0_esl_encoder_1_s0_writedata;                 // mm_interconnect_0:esl_encoder_1_s0_writedata -> esl_encoder_1:slave_writedata
	wire   [7:0] mm_interconnect_0_esl_encoder_1_s0_address;                   // mm_interconnect_0:esl_encoder_1_s0_address -> esl_encoder_1:slave_address
	wire         mm_interconnect_0_esl_encoder_1_s0_write;                     // mm_interconnect_0:esl_encoder_1_s0_write -> esl_encoder_1:slave_write
	wire         mm_interconnect_0_esl_encoder_1_s0_read;                      // mm_interconnect_0:esl_encoder_1_s0_read -> esl_encoder_1:slave_read
	wire  [31:0] mm_interconnect_0_esl_encoder_1_s0_readdata;                  // esl_encoder_1:slave_readdata -> mm_interconnect_0:esl_encoder_1_s0_readdata
	wire   [3:0] mm_interconnect_0_esl_encoder_1_s0_byteenable;                // mm_interconnect_0:esl_encoder_1_s0_byteenable -> esl_encoder_1:slave_byteenable
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // uart_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [esl_encoder_0:reset, esl_encoder_1:reset, esl_pwm_0:reset, esl_pwm_1:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sysid_qsys_0:reset_n, timer_0:reset_n, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	nios_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                             //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	nios_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	nios_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	nios_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.dataavailable (),                                          //                    .dataavailable
		.readyfordata  (),                                          //                    .readyfordata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	encoder_avalon_bus #(
		.DATA_WIDTH (32),
		.LED_WIDTH  (8)
	) esl_encoder_0 (
		.clk              (clk_clk),                                       //         clock_reset.clk
		.reset            (rst_controller_reset_out_reset),                //   clock_reset_reset.reset
		.slave_address    (mm_interconnect_0_esl_encoder_0_s0_address),    //                  s0.address
		.slave_read       (mm_interconnect_0_esl_encoder_0_s0_read),       //                    .read
		.slave_write      (mm_interconnect_0_esl_encoder_0_s0_write),      //                    .write
		.slave_readdata   (mm_interconnect_0_esl_encoder_0_s0_readdata),   //                    .readdata
		.slave_writedata  (mm_interconnect_0_esl_encoder_0_s0_writedata),  //                    .writedata
		.slave_byteenable (mm_interconnect_0_esl_encoder_0_s0_byteenable), //                    .byteenable
		.leds             (enc1leds_leds),                                 //      leds_interface.leds
		.encoder_a        (enc1a_encoder_a),                               // encoder_a_interface.encoder_a
		.encoder_b        (enc1b_encoder_b)                                // encoder_b_interface.encoder_b
	);

	encoder_avalon_bus #(
		.DATA_WIDTH (32),
		.LED_WIDTH  (8)
	) esl_encoder_1 (
		.clk              (clk_clk),                                       //         clock_reset.clk
		.reset            (rst_controller_reset_out_reset),                //   clock_reset_reset.reset
		.slave_address    (mm_interconnect_0_esl_encoder_1_s0_address),    //                  s0.address
		.slave_read       (mm_interconnect_0_esl_encoder_1_s0_read),       //                    .read
		.slave_write      (mm_interconnect_0_esl_encoder_1_s0_write),      //                    .write
		.slave_readdata   (mm_interconnect_0_esl_encoder_1_s0_readdata),   //                    .readdata
		.slave_writedata  (mm_interconnect_0_esl_encoder_1_s0_writedata),  //                    .writedata
		.slave_byteenable (mm_interconnect_0_esl_encoder_1_s0_byteenable), //                    .byteenable
		.leds             (enc2leds_leds),                                 //      leds_interface.leds
		.encoder_a        (enc2a_encoder_a),                               // encoder_a_interface.encoder_a
		.encoder_b        (enc2b_encoder_b)                                // encoder_b_interface.encoder_b
	);

	pwm_avalon_bus #(
		.DATA_WIDTH (32)
	) esl_pwm_0 (
		.clk              (clk_clk),                                   //       clock_reset.clk
		.reset            (rst_controller_reset_out_reset),            // clock_reset_reset.reset
		.slave_address    (mm_interconnect_0_esl_pwm_0_s0_address),    //                s0.address
		.slave_read       (mm_interconnect_0_esl_pwm_0_s0_read),       //                  .read
		.slave_write      (mm_interconnect_0_esl_pwm_0_s0_write),      //                  .write
		.slave_readdata   (mm_interconnect_0_esl_pwm_0_s0_readdata),   //                  .readdata
		.slave_writedata  (mm_interconnect_0_esl_pwm_0_s0_writedata),  //                  .writedata
		.slave_byteenable (mm_interconnect_0_esl_pwm_0_s0_byteenable), //                  .byteenable
		.ina              (pwma_ina),                                  //     pwm_interface.ina
		.inb              (pwma_inb),                                  //                  .inb
		.inc              (pwma_inc)                                   //                  .inc
	);

	pwm_avalon_bus #(
		.DATA_WIDTH (32)
	) esl_pwm_1 (
		.clk              (clk_clk),                                   //       clock_reset.clk
		.reset            (rst_controller_reset_out_reset),            // clock_reset_reset.reset
		.slave_address    (mm_interconnect_0_esl_pwm_1_s0_address),    //                s0.address
		.slave_read       (mm_interconnect_0_esl_pwm_1_s0_read),       //                  .read
		.slave_write      (mm_interconnect_0_esl_pwm_1_s0_write),      //                  .write
		.slave_readdata   (mm_interconnect_0_esl_pwm_1_s0_readdata),   //                  .readdata
		.slave_writedata  (mm_interconnect_0_esl_pwm_1_s0_writedata),  //                  .writedata
		.slave_byteenable (mm_interconnect_0_esl_pwm_1_s0_byteenable), //                  .byteenable
		.ina              (pwmb_ina),                                  //     pwm_interface.ina
		.inb              (pwmb_inb),                                  //                  .inb
		.inc              (pwmb_inc)                                   //                  .inc
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.nios2_qsys_0_instruction_master_readdatavalid    (nios2_qsys_0_instruction_master_readdatavalid),                //                                           .readdatavalid
		.esl_encoder_0_s0_address                         (mm_interconnect_0_esl_encoder_0_s0_address),                   //                           esl_encoder_0_s0.address
		.esl_encoder_0_s0_write                           (mm_interconnect_0_esl_encoder_0_s0_write),                     //                                           .write
		.esl_encoder_0_s0_read                            (mm_interconnect_0_esl_encoder_0_s0_read),                      //                                           .read
		.esl_encoder_0_s0_readdata                        (mm_interconnect_0_esl_encoder_0_s0_readdata),                  //                                           .readdata
		.esl_encoder_0_s0_writedata                       (mm_interconnect_0_esl_encoder_0_s0_writedata),                 //                                           .writedata
		.esl_encoder_0_s0_byteenable                      (mm_interconnect_0_esl_encoder_0_s0_byteenable),                //                                           .byteenable
		.esl_encoder_1_s0_address                         (mm_interconnect_0_esl_encoder_1_s0_address),                   //                           esl_encoder_1_s0.address
		.esl_encoder_1_s0_write                           (mm_interconnect_0_esl_encoder_1_s0_write),                     //                                           .write
		.esl_encoder_1_s0_read                            (mm_interconnect_0_esl_encoder_1_s0_read),                      //                                           .read
		.esl_encoder_1_s0_readdata                        (mm_interconnect_0_esl_encoder_1_s0_readdata),                  //                                           .readdata
		.esl_encoder_1_s0_writedata                       (mm_interconnect_0_esl_encoder_1_s0_writedata),                 //                                           .writedata
		.esl_encoder_1_s0_byteenable                      (mm_interconnect_0_esl_encoder_1_s0_byteenable),                //                                           .byteenable
		.esl_pwm_0_s0_address                             (mm_interconnect_0_esl_pwm_0_s0_address),                       //                               esl_pwm_0_s0.address
		.esl_pwm_0_s0_write                               (mm_interconnect_0_esl_pwm_0_s0_write),                         //                                           .write
		.esl_pwm_0_s0_read                                (mm_interconnect_0_esl_pwm_0_s0_read),                          //                                           .read
		.esl_pwm_0_s0_readdata                            (mm_interconnect_0_esl_pwm_0_s0_readdata),                      //                                           .readdata
		.esl_pwm_0_s0_writedata                           (mm_interconnect_0_esl_pwm_0_s0_writedata),                     //                                           .writedata
		.esl_pwm_0_s0_byteenable                          (mm_interconnect_0_esl_pwm_0_s0_byteenable),                    //                                           .byteenable
		.esl_pwm_1_s0_address                             (mm_interconnect_0_esl_pwm_1_s0_address),                       //                               esl_pwm_1_s0.address
		.esl_pwm_1_s0_write                               (mm_interconnect_0_esl_pwm_1_s0_write),                         //                                           .write
		.esl_pwm_1_s0_read                                (mm_interconnect_0_esl_pwm_1_s0_read),                          //                                           .read
		.esl_pwm_1_s0_readdata                            (mm_interconnect_0_esl_pwm_1_s0_readdata),                      //                                           .readdata
		.esl_pwm_1_s0_writedata                           (mm_interconnect_0_esl_pwm_1_s0_writedata),                     //                                           .writedata
		.esl_pwm_1_s0_byteenable                          (mm_interconnect_0_esl_pwm_1_s0_byteenable),                    //                                           .byteenable
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                           .clken
		.sysid_qsys_0_control_slave_address               (mm_interconnect_0_sysid_qsys_0_control_slave_address),         //                 sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata              (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),        //                                           .readdata
		.timer_0_s1_address                               (mm_interconnect_0_timer_0_s1_address),                         //                                 timer_0_s1.address
		.timer_0_s1_write                                 (mm_interconnect_0_timer_0_s1_write),                           //                                           .write
		.timer_0_s1_readdata                              (mm_interconnect_0_timer_0_s1_readdata),                        //                                           .readdata
		.timer_0_s1_writedata                             (mm_interconnect_0_timer_0_s1_writedata),                       //                                           .writedata
		.timer_0_s1_chipselect                            (mm_interconnect_0_timer_0_s1_chipselect),                      //                                           .chipselect
		.uart_0_s1_address                                (mm_interconnect_0_uart_0_s1_address),                          //                                  uart_0_s1.address
		.uart_0_s1_write                                  (mm_interconnect_0_uart_0_s1_write),                            //                                           .write
		.uart_0_s1_read                                   (mm_interconnect_0_uart_0_s1_read),                             //                                           .read
		.uart_0_s1_readdata                               (mm_interconnect_0_uart_0_s1_readdata),                         //                                           .readdata
		.uart_0_s1_writedata                              (mm_interconnect_0_uart_0_s1_writedata),                        //                                           .writedata
		.uart_0_s1_begintransfer                          (mm_interconnect_0_uart_0_s1_begintransfer),                    //                                           .begintransfer
		.uart_0_s1_chipselect                             (mm_interconnect_0_uart_0_s1_chipselect)                        //                                           .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
